module ex_5_32;
    reg A, B, C, D, E, F;
    reg A1, B1, C1, D1, E1, F1;

    initial 
    begin
        A = 1; B = 0; C = 0; D = 0; E = 1; F = 1;
    end

endmodule